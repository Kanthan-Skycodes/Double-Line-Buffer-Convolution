module cnn_first_layer#(
parameter imgDepth = 2,
parameter depth = 6,
parameter imgSize = 36,
parameter BUFFER_DEPTH = 256,
parameter DATA_WIDTH = 8,
parameter CHUNK_SIZE = 36,
parameter NUM_PORTS = 2,
parameter DEPTH = CHUNK_SIZE * NUM_PORTS * 4, // larger for multiple chunks
parameter ADDR_WIDTH = 9
)(
input clk,
input rst,
output signed [42:0] maxpool_out,
output signed [25:0] relu_out_1,
output done_o1,
output control
);
// Interconnecting signals
wire signed [25:0] dout0;
wire signed [25:0] out_1;
wire wr_en;
wire signed [42:0]result;
wire done;
// Control signals generated by the FSM
reg done_i1;
reg start1;
reg rd_en;
// FSM state definition
reg [3:0] state;
localparam
S0 = 0, // Wait after reset (2 cycles)
S1 = 1, // Assert start1 pulse (one cycle)
S11 = 8,
S2 = 2, // Wait 57 cycles for first-layer phase (done_i1/wr_en active)
S3 = 3, // End first-layer phase (deassert done_i1/wr_en)
S4 = 4, // Assert start2 pulse (one cycle)
S41 = 9,
S42 = 10,
S43 = 11,
S5 = 5, // Wait 57 cycles for second-layer phase (done_i2 and rd_en active)
S6 = 6, // End second-layer phase (deassert done_i2 and rd_en)
S_IDLE= 7; // Idle/finish state
// Counter signals and reset control
reg [31:0] counter;
reg counter_reset;
assign wr_en = done_i1 && done_o1;
//-------------------------------------------------------------------------
// Instantiate the First Layer module
//-------------------------------------------------------------------------
first_layer#(imgDepth, depth, imgSize) firstLayer (
.clk(clk),
.rst(rst),
.done_i(done_i1),
.start(start1),
.out(relu_out_1),
.done_o(done_o1)
);
/////////////////////////////////////////////
//////relu
//////////////////////////////////////////////
relu r1(
.in(out_1),
.out()
);

///////////////////////////////////////////////////////////////////////////
// maxpool block
//////////////////////////////////////////////////////////////////////////
top_for_maxpool max(
.d_in(relu_out_1),
.clk(clk),
.rst(rst),
.done_i(done_o1),
.max(maxpool_out),
.done_o(done),
.control(control)
);
//-------------------------------------------------------------------------
// COUNTER BLOCK (Runs Independently)
//-------------------------------------------------------------------------
always @(posedge clk) begin
if (rst)
counter <= 0;
else if (counter_reset)
counter <= 0;
else
counter <= counter + 1;
end
//-------------------------------------------------------------------------
// FSM BLOCK: State transitions and control signal assignments.
// Notice we have separated the pulse states (S1 and S4) from the waiting states.
//-------------------------------------------------------------------------
always @(posedge clk) begin
if (rst) begin
state <= S0;
start1 <= 0;
start2 <= 0;
rd_en <= 0;
done_i1 <= 0;
done_i2 <= 0;
counter_reset <= 1; // Reset counter immediately after reset.
end else begin
// By default, deassert counter_reset.
counter_reset <= 0;
case (state)
S0: begin
// Wait for 2 cycles after reset
if (counter >= 2) begin
state <= S1;
counter_reset <= 1; // Reset counter for next state timing.
end
end
S1: begin
// Assert start1 for one full clock cycle.
start1 <= 1;
// Transition in the next clock cycle.
state <= S11;
counter_reset <= 1; // Reset counter to start 57-cycle count.
end
S11:begin
state <= S2;
end
S2: begin
// Deassert start1 (pulse ended) and drive done_i1.
start1 <= 0;
done_i1 <= 1;
// Drive wr_en conditionally on done_o1.
if (counter >= 1370+(imgSize*imgDepth)) begin
state <= S3;
counter_reset <= 1;
end
end
S3: begin
// Deassert done_i1 and wr_en, then move to second phase.
done_i1 <= 0;
state <= S_IDLE;
end

S_IDLE: begin
// Idle state; no further transitions.
end
default: state <= S_IDLE;
endcase
end
end
endmodule

module first_layer#(parameter imgDepth=2,parameter depth=5,parameter imgSize=25)(
input clk,
input rst,
input done_i,
input start,
output signed [25:0]out,
output done_o
);
wire signed [8:0]in;
localparam path="testKernelWeights.txt";
image_provider #(imgSize,imgDepth) prov(
.clk(clk),
.rst(rst),
.start(start),
.pixel_data(in),
.pixel_valid()
);
processElement#(imgDepth,depth,path) pe(
.clk(clk),
.rst(rst),
.grayscale_i(in),
.done_i(done_i),
.out(out),
.done_o(done_o)
);
endmodule
/////////////////////////////////////////////image_provider/////////////////////////////////////////////
module image_provider #(parameter imgSize = 36, parameter imgDepth = 1)(
input clk,
input rst,
input start,
output reg signed [8:0] pixel_data,
output reg pixel_valid
);
reg signed [8:0] rom [0:imgSize-1]; // ROM to store image data
reg [31:0] addr; // Address pointer for ROM
reg [31:0] depth_counter; // Counter for imgDepth
reg [1:0] state; // FSM state
// Initialize ROM with image data
initial begin
$readmemb("camera_binary.txt", rom); // Load image data from file
end
// FSM to control image data read
always @(posedge clk or posedge rst) begin
if (rst) begin
state <= 0;
addr <= 0;
depth_counter <= 0;
pixel_data <= 0;
pixel_valid <= 0;
end else begin
case (state)
0: begin // Idle state
if (start) begin
state <= 1;
addr <= 0;
depth_counter <= 0;
pixel_valid <= 1;
end
end
1: begin // Read and output pixel data continuously
pixel_data <= rom[addr];
if (addr < imgSize - 1) begin
addr <= addr + 1;
end else if (depth_counter < imgDepth - 1) begin
depth_counter <= depth_counter + 1;
addr <= 0; // Restart image output without gap
end else begin
state <= 0;
pixel_valid <= 0;
end
end
endcase
end
end
endmodule
//////////////////////////////////////////////////processing Element for first layer(ch)////////////////////////////////////////
module processElement#(parameter imgDepth=64,parameter depth=128,parameter
path="testKernelWeights.txt" )(
input clk,
input rst,
input signed [8:0]grayscale_i,
input done_i,
output signed [25:0]out,
output done_o
);
wire signed [8:0]w0,w1,w2,w3,w4,w5,w6,w7,w8;
imageControl#(imgDepth,depth) imgC(
.clk(clk),
.rst(rst),
.grayscale_i(grayscale_i),
.done_i(done_i),
// .ut [24:0]conv_out,
.d0_o(w0),
.d1_o(w1),
.d2_o(w2),
.d3_o(w3),
.d4_o(w4),
.d5_o(w5),
.d6_o(w6),
.d7_o(w7),
.d8_o(w8),
.done_o(done_o));
conv_top#(imgDepth,path) ct
(
.clk(clk),
.rst(rst),
.in0(w0),
.in1(w1),
.in2(w2),
.in3(w3),
.in4(w4),
.in5(w5),
.in6(w6),
.in7(w7),
.in8(w8),
.done_o(done_o),//
.out(out)
);
endmodule
module imageControl#(parameter imgDepth=2,parameter depth=5)(
input clk,
input rst,
input signed [8:0] grayscale_i,
input done_i,
// output [24:0]conv_out,
output signed [8:0] d0_o,
output signed [8:0] d1_o,
output signed [8:0] d2_o,
output signed [8:0] d3_o,
output signed [8:0] d4_o,
output signed [8:0] d5_o,
output signed [8:0] d6_o,
output signed [8:0] d7_o,
output signed [8:0] d8_o,
output done_o
);
wire signed [8:0] double_line_fifo_data0;
wire signed [8:0] double_line_fifo_data1;
wire signed [8:0] double_line_fifo_data2;
wire double_line_fifo_done;
doubleLineBuffer #(depth)db (
.clk(clk),
.rst(rst),
.we(done_i),
.data_i(grayscale_i),
.data0_o(double_line_fifo_data0),
.data1_o(double_line_fifo_data1),
.data2_o(double_line_fifo_data2),
.done_o(double_line_fifo_done)
);
striding #(imgDepth,depth)SD(
.clk(clk),
.rst(rst),
.d0_i(double_line_fifo_data0),
.d1_i(double_line_fifo_data1),
.d2_i(double_line_fifo_data2),
.done_i(double_line_fifo_done),
.d0_o(d0_o),
.d1_o(d1_o),
.d2_o(d2_o),
.d3_o(d3_o),
.d4_o(d4_o),
.d5_o(d5_o),
.d6_o(d6_o),
.d7_o(d7_o),
.d8_o(d8_o),
.done_o(done_o)
);
endmodule
////////////////////////////////////double Line Buffer Module(ch)///////////////////////////////////////
module doubleLineBuffer#(parameter depth=5)(
input clk,
input rst,
input we,
input signed[8:0]data_i,
output signed [8:0]data0_o,
output signed [8:0]data1_o,
output signed [8:0]data2_o,
output done_o
);
wire signed [8:0]fifo1;
wire signed [8:0]fifo2;
wire fifo1_done,fifo2_done;
assign data0_o = data_i;
assign data1_o = fifo1;
assign data2_o = fifo2;
assign done_o = fifo1_done;
lineBuffer #(depth) lbo (
.clk(clk),
.rst(rst),
. we(we),
.data_i(data_i),
.data_o(fifo1),
. done_o(fifo1_done)
);
lineBuffer #(depth)lb1 (
.clk(clk),
.rst(rst),
.we(fifo1_done),
.data_i(fifo1),
.data_o(fifo2),
.done_o(fifo2_done)
);
endmodule
//////////////////////////////////////////Line Buffer Module(ch)/////////////////////////////////////////////
module lineBuffer#(parameter depth=5)(
input clk,
input rst,
input we,
input signed [8:0] data_i,
// input done_i,
output signed [8:0] data_o,
output done_o
);
// parameter depth = 640;
//for normal checking we can use this
reg signed [25:0] mem [0:depth-1];
reg [9:0] rd_pointer; ///////////////image is 240x240 then 240 we will get with 8 bits////////
reg [9:0] wr_pointer;
reg [9:0] i_counter;
assign done_o = (i_counter == depth) ? 1:0;
assign data_o = mem[rd_pointer];
/////////////////////////////counting the pixel /////////
always@(posedge clk)
begin
if(rst)
begin
i_counter<=0;
end
else
begin
if(we == 1)
begin
i_counter <= (i_counter == depth) ? i_counter:i_counter+1;
end
end
end
////////////////////////////writing////////////////
always@(posedge clk)
begin
if(rst)
begin
wr_pointer<= 0;
end
else
begin
if( we==1)
begin
mem[wr_pointer] <= data_i;
wr_pointer <= (wr_pointer == depth-1)? 0: wr_pointer+1;
end
end
end
//////////////////////////////////reading///////////////////////
always@(posedge clk)
begin
if(rst)
begin
rd_pointer <= 0;
end
else
begin
if( we==1)
begin
if(i_counter == depth)
begin
rd_pointer <= (rd_pointer == depth-1) ? 0: rd_pointer+1;
end
end
end
end
endmodule
//////////////////////////////////////////////////////////Striding Module(ch
important)/////////////////////////////////////////////////////////
`define imgSize 512*512
module striding#(parameter imgDepth=2, parameter depth=4)(
input clk,
input rst,
input signed[8:0]d0_i,
input signed[8:0]d1_i,
input signed[8:0]d2_i,
input done_i,
output reg signed [8:0] d0_o,d1_o,d2_o,d3_o,d4_o,d5_o,d6_o,d7_o,d8_o,
output done_o
);
localparam row= depth;
localparam col= depth;
reg [8:0] data0,data1,data2,data3,data4,data5,data6,data7,data8;
reg [7:0] i_counter;
reg [9:0] irow,icol;
assign done_o = (i_counter==2)?1:0;
always@(posedge clk)
begin
if(rst)
begin
irow <= 0;
icol <= 0;
end
else
begin
if(done_o == 1)
begin
icol <= (icol == col-1)?0:icol+1;
if(icol == col-1)
irow <= (irow == row-1)?0:irow+1;
end
end
end
always@(*)
begin
if(rst)
begin
d0_o<=0;
d1_o<=0;
d2_o<=0;
d3_o<=0;
d4_o<=0;
d5_o<=0;
d6_o<=0;
d7_o<=0;
d8_o<=0;
end
else
begin
if(done_o == 1)
begin
////////////pos1/////////////
if(irow ==0 && icol ==0)
begin
d0_o<=0;
d1_o<=0;
d2_o<=0;
d3_o<=0;
d4_o<=data4;
d5_o<=data5;
d6_o<=0;
d7_o<=data7;
d8_o<=data8;
end
//////////////////////pos2///////////
else
if(irow == 0 && icol > 0 && icol < col-1)
begin
d0_o<=0;
d1_o<=0;
d2_o<=0;
d3_o<=data3;
d4_o<=data4;
d5_o<=data5;
d6_o<=data6;
d7_o<=data7;
d8_o<=data8;
end
///////////////////pos3////////////
else
if(irow == 0 && icol == col-1)
begin
d0_o<=0;
d1_o<=0;
d2_o<=0;
d3_o<=data3;
d4_o<=data4;
d5_o<=0;
d6_o<=data6;
d7_o<=data7;
d8_o<=0;
end
/////////////////////////pos4/////////////////////////
else
if(irow > 0 && irow < row-1 && icol == 0)
begin
d0_o<=0;
d1_o<=data1;
d2_o<=data2;
d3_o<=0;
d4_o<=data4;
d5_o<=data5;
d6_o<=0;
d7_o<=data7;
d8_o<=data8;
end
///////////////////////////////pos5////////////////
else
if (irow > 0 && irow < row-1 && icol > 0 && icol < col-1)
begin
d0_o<=data0;
d1_o<=data1;
d2_o<=data2;
d3_o<=data3;
d4_o<=data4;
d5_o<=data5;
d6_o<=data6;
d7_o<=data7;
d8_o<=data8;
end
///////////////////////////////////////pos6//////////////////
else
if(irow > 0 && irow < row-1 && icol == col-1)
begin
d0_o<=data0;
d1_o<=data1;
d2_o<=0;
d3_o<=data3;
d4_o<=data4;
d5_o<=0;
d6_o<=data6;
d7_o<=data7;
d8_o<=0;
end
////////////////////////////pos7/////////////////////
else
if(irow == row-1 && icol == 0)
begin
d0_o<=0;
d1_o<=data1;
d2_o<=data2;
d3_o<=0;
d4_o<=data4;
d5_o<=data5;
d6_o<=0;
d7_o<=0;
d8_o<=0;
end
///////////////////////////pos8////////////////////////////
else
if(irow == row-1 && icol > 0 && icol < col-1)
begin
d0_o<=data0;
d1_o<=data1;
d2_o<=data2;
d3_o<=data3;
d4_o<=data4;
d5_o<=data5;
d6_o<=0;
d7_o<=0;
d8_o<=0;
end
//////////////////////////pos9///////////////////
else
if ( irow == row-1 && icol == col-1)
begin
d0_o<=data0;
d1_o<=data1;
d2_o<=0;
d3_o<=data3;
d4_o<=data4;
d5_o<=0;
d6_o<=0;
d7_o<=0;
d8_o<=0;
end
end
end
end
always@(posedge clk)
begin
if(rst)
begin
i_counter<=0;
end
else
begin
if(done_i==1)
begin
i_counter<=(i_counter == 2)? i_counter:i_counter+1;
end
end
end
always@(posedge clk)
begin
if(rst)
begin
data0<=0;
data1<=0;
data2<=0;
data3<=0;
data4<=0;
data5<=0;
data6<=0;
data7<=0;
data8<=0;
end
else
begin
if(done_i==1)
begin
data0<=data1;
data1<=data2;
data2<=d2_i;
data3<=data4;
data4<=data5;
data5<=d1_i;
data6<=data7;
data7<=data8;
data8<=d0_i;
end
end
end
endmodule
///////////////////////////////////////////////////////////multiply and accumulate /////////////////////////////////////////////
module conv_top#(parameter imgDepth = 2,parameter
path="testKernelWeights.txt")(clk,rst,in0,in1,in2,in3,in4,in5,in6,in7,in8,done_o,out);
input clk,rst;
input signed [8:0]in0,in1,in2,in3,in4,in5,in6,in7,in8;
input done_o;
output signed [25:0]out;
wire signed [8:0]k0,k1,k2,k3,k4,k5,k6,k7,k8;
wire signed [25:0]res;
krom11#(imgDepth,path) rom(
.clk(clk),
.rst(rst),
.data0(k0),
.data1(k1),
.data2(k2),
.data3(k3),
.data4(k4),
.data5(k5),
.data6(k6),
.data7(k7),
.data8(k8)
);
convolution c0(
.clk(clk),
.rst(rst),
.in0(in0),
.in1(in1),
.in2(in2),
.in3(in3),
.in4(in4),
.in5(in5),
.in6(in6),
.in7(in7),
.in8(in8),
.b0(k0),
.b1(k1),
.b2(k2),
.b3(k3),
.b4(k4),
.b5(k5),
.b6(k6),
.b7(k7),
.b8(k8),
.conv_out(out));
endmodule
module convolution
(clk,rst,in0,in1,in2,in3,in4,in5,in6,in7,in8,b0,b1,b2,b3,b4,b5,b6,b7,b8,conv_out);
input signed [8:0]in0,in1,in2,in3,in4,in5,in6,in7,in8;
input signed [8:0]b0,b1,b2,b3,b4,b5,b6,b7,b8;
input clk,rst;
output signed [25:0]conv_out;
wire signed [16:0]mul0,mul1,mul2,mul3,mul4,mul5,mul6,mul7,mul8;
wire signed [24:0]sum_out_int,sum_out;
multiply m0(in0,b0,mul0);
multiply m1(in1,b1,mul1);
multiply m2(in2,b2,mul2);
multiply m3(in3,b3,mul3);
multiply m4(in4,b4,mul4);
multiply m5(in5,b5,mul5);
multiply m6(in6,b6,mul6);
multiply m7(in7,b7,mul7);
multiply m8(in8,b8,mul8);
assign conv_out = (mul0 + mul1 + mul2 + mul3 + mul4 + mul5 + mul6 + mul7 + mul8);
//assign conv_out = sum_out_int /9;//assign conv_out = sum_out_int /9;
//accumulator #(imgDepth)a0(.clk(clk),.rst(rst),.in(sum_out),.out(conv_out));
endmodule
//////////////////////////////////////////////////multiply module////////////////////////////////////////////////////
module multiply(
input signed [8:0]a,
input signed [8:0]b,
output reg signed [16:0]mul
);
always@(*)
begin
mul <= a*b;
end
endmodule
///////////////////////////////////////////relu for first layer////////////////////////////////////////////////////
module relu(
input [25:0]in,
output reg [25:0]out
);
always@(*)
begin
if(in[25] == 1'b1)
out <= 0;
else
out <= in;
end
endmodule
//////////////////////////////////////////////////Maxpool///////////////////////////////////////////////////////
module top_for_maxpool(
input [42:0]d_in,
input clk,
input rst,
input done_i,
output [42:0]max,
output done_o,
output control
);
wire [42:0]out;
wire en1,en2;
wire done_o2;
max_finder_for_elements
t2(.d_in(d_in),.clk(clk),.done_i(done_i),.rst(rst),.max_of_two(out),.enable_out(en1),.done_o(done
_o2));
max_finder_for_rows
t3(.d_in(out),.clk(clk),.rst(rst),.done_i(done_i),.d_out(max),.done_o(done_o),.en1(en2));
write_controller w1(.a(en1),.b(clk),.c(done_o),.d(en2),.control(control));
endmodule
///////////////////////////////////////maxfinder for elements//////////////////////////////////////////////////
module max_finder_for_elements(
input [42:0]d_in,
input clk,rst,
input done_i,
output [42:0]max_of_two,
output enable_out,
output done_o
);
wire [42:0]out;
reg [24:0]i_counter;
assign done_o = (i_counter == 2)?1:0;
en_gen_for_two_elements e1(.clk(clk),.rst(rst),.en(enable_out));
dflipflop d1(.d_in(d_in),.clk(clk),.rst(rst),.d_out(out));
max_finder_with_enable m1(.a(out),.b(d_in),.enable(~enable_out),.max(max_of_two));
always@(posedge clk)
begin
if(rst)
begin
i_counter<=0;
end
else
begin
if(done_i==1)
begin
i_counter<=(i_counter == 2)? i_counter:i_counter+1;
end
end
end
endmodule
///////////////////////////////////////////enable generator for two elements///////////////////////////////
module en_gen_for_two_elements(
input clk,
input rst,
output reg en
);
reg state = 1'b0;
always @(posedge clk or posedge rst) begin
if (rst) begin
state <= 1'b1;
en <= 1'b0; // Initialize enable to 0 on reset
end else begin
state <= ~state;
en <= state;
end
end
endmodule
////////////////////////////////////////////d flipflop//////////////////////////////////////////////////////
module dflipflop(
input [42:0]d_in,
input clk,
input rst,
output reg [42:0]d_out
);
reg [42:0]temp;
always@(posedge clk or posedge rst)
begin
if(rst) begin
temp <= 0;
d_out <= 0;
end
else
temp <= d_in;
end
always@(posedge clk)
begin
d_out <= temp;
end
endmodule
/////////////////////////////////////max finder for two elements///////////////////////////////////////
module max_finder_with_enable(
input [42:0]a,
input [42:0]b,
input enable,
output reg [42:0]max
);
always@(posedge enable)
begin
max <= (a>b) ? a : b;
end
endmodule
///////////////////////////////////max_finder for rows//////////////////////////////////////////////
module max_finder_for_rows(
input [42:0]d_in,
input clk,
input rst,
input done_i,
output [42:0]d_out,
output done_o,
output en1
);
wire [42:0]out;
freq_divider f1(.clk(clk),.rst(rst),.done_o(done_o),.n(32'd128),.enable(en1));
lineBuffer_for_max
lb1(.clk(clk),.rst(rst),.we(done_i),.data_i(d_in),.data_o(out),.done_o(done_o));
max_for_buffer m2(.a(d_in),.b(out),.start(done_o),.enable(en1),.max(d_out));
endmodule
/////////////////////////////////////frequency divider///////////////////////////////////////////
module freq_divider (
input wire clk, // Input clock of frequency f
input wire rst, // Reset signal
input wire done_o, // Signal from top module to start counting delay
input wire [31:0] n, // Divider factor n (frequency division factor)
output reg enable // Output enable signal with frequency f/n
);
reg [31:0] counter; // Single counter for delay and frequency division
reg enable_active; // Flag to switch from delay to frequency division
// Calculate half of n
wire [31:0] half_n = n >> 1;
always @(posedge clk or posedge rst) begin
if (rst) begin
counter <= 0; // Initialize counter
enable <= 0;
enable_active <= 0; // Disable enable output initially
end else if (!enable_active && done_o) begin
// Delay phase: wait for n/2 clock cycles after done_o is high
if (counter == (half_n - 1)) begin
enable_active <= 1; // Activate enable after n/2 clock pulses
counter <= 0; // Reset counter for frequency division
enable <= 1; // Set enable high immediately after delay
end else begin
counter <= counter + 1;
end
end else if (enable_active) begin
// Frequency division phase
if (counter == (n - 1)) begin
counter <= 0;
enable <= ~enable; // Toggle enable every n clock cycles
end else begin
counter <= counter + 1;
end
end
end
endmodule
//////////////////////////////////////////////////line buffer////////////////////////////////////////////////////
module lineBuffer_for_max(
input clk,
input rst,
input we,
input [42:0] data_i,
// input done_i,
output [42:0] data_o,
output done_o
);
// parameter depth = 640;
parameter depth = 128; //for normal checking we can use this
reg [42:0] mem [0:depth-1];
reg [9:0] rd_pointer; ///////////////image is 240x240 then 240 we will get with 8 bits////////
reg [9:0] wr_pointer;
reg [9:0] i_counter;
assign done_o = (i_counter == depth) ? 1:0;
assign data_o = mem[rd_pointer];
/////////////////////////////counting the pixel /////////
always@(posedge clk)
begin
if(rst)
begin
i_counter<=0;
end
else
begin
if(we == 1)
begin
i_counter <= (i_counter == depth) ? i_counter:i_counter+1;
end
end
end
////////////////////////////writing////////////////
always@(posedge clk)
begin
if(rst)
begin
wr_pointer<= 0;
end
else
begin
if( we==1)
begin
mem[wr_pointer]<= data_i;
wr_pointer <= ( wr_pointer ==depth-1)? 0: wr_pointer+1;
end
end
end
//////////////////////////////////reading///////////////////////
always@(posedge clk)
begin
if(rst)
begin
rd_pointer <= 0;
end
else
begin
if( we==1)
begin
if(i_counter == depth)
begin
rd_pointer <= (rd_pointer == depth-1) ? 0: rd_pointer+1;
end
end
end
end
endmodule
////////////////////////////////////////////////////////////////max for two elements in different rows/////////////////
module max_for_buffer(
input [42:0]a,
input [42:0]b,
input start,
input enable,
output reg [42:0]max
);
always@(*)
begin
if(start && enable)
begin
max <= (a>b)?a:b;
end
end
endmodule
